module bridge_design();

endmodule
